library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity i2s_loop_tb is

end entity;

architecture arch of i2s_loop_tb is

begin

end architecture;
