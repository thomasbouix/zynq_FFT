library ieee;
use ieee.std_logic_1164.all;

entity vga_controller_tb is 

end entity;

architecture arc_vga_controller_tb of vga_controller_tb is

begin	

end arc_vga_controller_tb;

